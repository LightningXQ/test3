library verilog;
use verilog.vl_types.all;
entity TB_not_gate is
end TB_not_gate;
